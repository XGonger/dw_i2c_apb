//=======================================================================
// COPYRIGHT (C) 2018-2020 RockerIC, Ltd.
// This software and the associated documentation are confidential and
// proprietary to RockerIC, Ltd. Your use or disclosure of this software
// is subject to the terms and conditions of a consulting agreement
// between you, or your company, and RockerIC, Ltd. In the event of
// publications, the following notice is applicable:
//
// ALL RIGHTS RESERVED
//
// The entire notice above must be reproduced on all authorized copies.
//
// VisitUs  : www.rockeric.com
// Support  : support@rockeric.com
// WeChat   : eva_bill 
//-----------------------------------------------------------------------
`ifndef LVC_I2C_MASTER_DRIVER_COMMON_SV
`define LVC_I2C_MASTER_DRIVER_COMMON_SV

class lvc_i2c_master_driver_common extends lvc_i2c_bfm_common;

  `uvm_object_utils_begin(lvc_i2c_master_driver_common)
  `uvm_object_utils_end
  semaphore      lock;            //if current send the restart cmd, next transaction need not to send start cmd
  bit            nack_flag=0;     // flag about nack generated by slave
  bit is10bits_again=0;
  bit same_slv_addr_in10bit=0;
  bit [9:0] pre_addr=0;
  extern function new(string name = "lvc_i2c_master_driver_common");

  extern virtual task send_xact(lvc_i2c_master_transaction trans);
  extern virtual task collect_response_from_vif(lvc_i2c_master_transaction trans);
  extern task start_gen();
  extern task stop_gen();
  extern task rw_slave_7bit_addr(bit[6:0] addr, bit rw);
  extern task rw_slave_10bit_addr(bit [9:0] addr, bit rw);
  extern task send_byte(bit[7:0] send_byte);
  extern task recv_byte(output bit[7:0] recv_data);
  extern task recv_byte_noack(output bit[7:0] recv_data);
  extern task send_start_byte();
  extern task pre_hs_in_fm_send_byte(bit[7:0] send_byte);
  extern task pre_hs_in_fm_plus_send_byte(bit[7:0] send_byte);
  extern task pre_hs_in_fm_start_gen();
  extern task pre_hs_in_fm_plus_start_gen();
  extern task re_start_gen();
  extern task drive_data(lvc_i2c_master_transaction trans);
  extern task rw_same_slave_10bit_addr(bit [9:0] addr, bit rw);

endclass

function lvc_i2c_master_driver_common::new(string name = "lvc_i2c_master_driver_common");
  super.new(name);
  lock = new(1);
endfunction

task lvc_i2c_master_driver_common::send_xact(lvc_i2c_master_transaction trans);
  lvc_i2c_master_transaction trans_temp;
    clk_low_offset_gen();
    drive_data(trans);
endtask

task lvc_i2c_master_driver_common::drive_data(lvc_i2c_master_transaction trans);
  bit       rw;   //0--write, 1--read
  bit[7:0]  recv_data;
  bit[7:0]  gen_call_first_byte = 8'b0000_0000;
  bit[7:0]  gen_call_second_byte = trans.sec_byte_gen_call;
  bit[7:0]  device_id_w = 8'b1111_1000;
  bit[7:0]  device_id_r = 8'b1111_1001;
  bit[7:0]  hs_code     = {5'b00001,cfg.master_code};
  bit[2:0]  num_of_retry=0;

  if(trans.retry_if_nack) 
      num_of_retry = trans.num_of_retry;
  else
      num_of_retry=0;

  case(trans.cmd)
    I2C_WRITE:
      for(int retry_num=0; retry_num<=num_of_retry; ) begin
          nack_flag = 0;
          if(cfg.bus_speed == HIGHSPEED_MODE) begin
              if(cfg.start_hs_in_fm_plus==0) begin
                  pre_hs_in_fm_start_gen();
                  pre_hs_in_fm_send_byte(hs_code);
              end else begin
                  pre_hs_in_fm_plus_start_gen();
                  pre_hs_in_fm_plus_send_byte(hs_code);
              end

              re_start_gen();

              if(trans.addr_10bit ==1)
                  rw_slave_10bit_addr(trans.addr, 0);
              else
                  rw_slave_7bit_addr(trans.addr[6:0], 0);

              // check and response when addr/send_start_byte nack generated by slave    
              if(nack_flag==1) begin
                  if(num_of_retry==0 | !trans.retry_if_nack) begin
                      stop_gen();
                      return;
                  end
                  else if(retry_num==num_of_retry) begin
                      retry_num++; 
                      continue;
                  end
                  else begin
                      retry_num++;
                      if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                          stop_gen();
                      else
                          re_start_gen();
                      continue;
                  end
              end  //if(nack_flag==1)
            
              for(int i=0; i<trans.data.size();i++)
              begin
                  send_byte(trans.data[i]);
                  // check and response when data nack generated by slave    
                  if(nack_flag==1) begin
                      if(num_of_retry==0 | !trans.retry_if_nack) begin
                          stop_gen();
                          return;
                      end
                      else if(retry_num==num_of_retry) begin
                          retry_num++;
                          continue;
                      end
                      else begin
                          retry_num++;
                          if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                              stop_gen();
                          else
                              re_start_gen();
                          break;
                      end
                  end //if(nack_flag==1)
              end//for(int i=0; i<trans.data.size();i++)
              
              if(nack_flag==0 | retry_num==num_of_retry+1) begin
                  if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                      stop_gen();
                  else
                      re_start_gen();
                  break;
              end //if(nack_flag==0)
          end //if(cfg.bus_speed == HIGHSPEED_MODE)
          else begin
              start_gen();
            
              if(trans.send_start_byte == 1)
                  send_start_byte();
           
              if(trans.addr_10bit ==1) begin
                  is10bits_again=1;
                  pre_addr=trans.addr;

                  rw_slave_10bit_addr(trans.addr, 0);
              end else
                  rw_slave_7bit_addr(trans.addr[6:0], 0);
            
              // check and response when addr/send_byte nack generated by slave    
              if(nack_flag==1) begin
                  if(num_of_retry==0 | !trans.retry_if_nack) begin
                      stop_gen();
                      return;
                  end
                  else if(retry_num==num_of_retry) begin
                      retry_num++;
                      continue;
                  end
                  else begin
                      retry_num++;
                      if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                          stop_gen();
                      else
                          re_start_gen();                      
                      continue;
                  end
                 // if(retry_num==trans.num_of_retry | !trans.retry_if_nack) begin
                 //     stop_gen();
                 //     return;
                 // end
                 // else begin
                 //     re_start_gen();
                 //     continue;
                 // end
              end //if(nack_flag==1)
            
              for(int i=0; i<trans.data.size();i++)
              begin
                  send_byte(trans.data[i]);
                  // check and response when data nack generated by slave    
                  if(nack_flag==1) begin
                      if(num_of_retry==0 | !trans.retry_if_nack) begin
                          stop_gen();
                          return;
                      end
                      else if(retry_num==num_of_retry) begin
                          retry_num++;
                          continue;
                      end
                      else begin
                          retry_num++;
                          if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                              stop_gen();
                          else
                              re_start_gen();
                          break;
                      end
                  end
              end  //for(int i=0; i<trans.data.size();i++)
            
              if(nack_flag==0 | retry_num==num_of_retry+1) begin
                  if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                      stop_gen();
                  else
                      re_start_gen();
                  break;
              end  //if(nack_flag==0)
          end  //else high_speed
      end //for(int i=0; i<=trans.num_of_retry; i++)
    I2C_READ: 
      for(int retry_num=0; retry_num<=num_of_retry; ) begin  
          if(cfg.bus_speed == HIGHSPEED_MODE) begin
              if(cfg.start_hs_in_fm_plus==0) begin//start hs in fm speed
                  pre_hs_in_fm_start_gen();
                  pre_hs_in_fm_send_byte(hs_code);
              end else begin
                  pre_hs_in_fm_plus_start_gen();
                  pre_hs_in_fm_plus_send_byte(hs_code);
              end
            
              re_start_gen();
            
              if(trans.addr_10bit ==1)
                  rw_slave_10bit_addr(trans.addr, 1);
              else
                  rw_slave_7bit_addr(trans.addr[6:0], 1);

              // check and response when addr/send_start_byte nack generated by slave    
              if(nack_flag==1) begin
                  if(num_of_retry==0 | !trans.retry_if_nack) begin
                      stop_gen();
                      return;
                  end
                  else if(retry_num==num_of_retry) begin
                      retry_num++; 
                      continue;
                  end
                  else begin
                      retry_num++;
                      if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                          stop_gen();
                      else
                          re_start_gen();
                      continue;
                  end
              end //if(nack_flag==1)

              for(int i=0; i<trans.data.size();i++)
              begin
                  recv_byte(recv_data);
                  trans.data[i] = recv_data;
              end
              //received last byte data and master send out nack to slave
              recv_byte_noack(recv_data);
              trans.data[trans.data.size()-1] = recv_data;
               
              if(trans.sr_or_p_gen==0  | retry_num==num_of_retry+1  | retry_num==0) begin //0--gen sotp, 1--gen re-start
                  retry_num++;
                  stop_gen();
              end
              else
                  re_start_gen();
          end  //if(cfg.bus_speed == HIGHSPEED_MODE)
          else begin
              start_gen();
            
              if(trans.send_start_byte == 1)
                  send_start_byte();
            
              if(trans.addr_10bit ==1) begin
                if(is10bits_again==0) begin
                  rw_slave_10bit_addr(trans.addr, 1);
                end else if(is10bits_again==1) begin
                  if(trans.addr==pre_addr) begin
                    rw_same_slave_10bit_addr(trans.addr, 1);
                  end else begin
                    rw_slave_10bit_addr(trans.addr, 1);
                  end
                end
              end else begin
                  rw_slave_7bit_addr(trans.addr[6:0], 1);
              end
              // check and response when addr/send_start_byte nack generated by slave    
              if(nack_flag==1) begin
                  if(num_of_retry==0 | !trans.retry_if_nack) begin
                      stop_gen();
                      return;
                  end
                  else if(retry_num==num_of_retry) begin
                      retry_num++; 
                      continue;
                  end
                  else begin
                      retry_num++;
                      if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                          stop_gen();
                      else
                          re_start_gen();
                      continue;
                  end
              end  //if(nack_flag==1)
            
              for(int i=0; i<trans.data.size()-1;i++)
                begin
                    recv_byte(recv_data);
                    trans.data[i] = recv_data;
                end
              recv_byte_noack(recv_data);
              trans.data[trans.data.size()-1] = recv_data;
            
              if(trans.sr_or_p_gen==0  | retry_num==num_of_retry+1  | retry_num==0) begin //0--gen sotp, 1--gen re-start
                  retry_num++;
                  stop_gen();
              end
              else
                  re_start_gen();              
          end  ///else
      end//for(int retry_num=0; retry_num<=trans.num_of_retry; )
    I2C_GEN_CALL: 
      for(int retry_num=0; retry_num<=num_of_retry;) begin  
          start_gen();
          
          if(trans.send_start_byte==1)
              send_start_byte();
          
          send_byte(gen_call_first_byte);
          // check and response when addr/send_start_byte nack generated by slave    
          if(nack_flag==1) begin
              if(num_of_retry==0 | !trans.retry_if_nack) begin
                  stop_gen();
                  return;
              end
              else if(retry_num==num_of_retry) begin
                  retry_num++;
                  continue;
              end
              else begin
                  retry_num++;
                  if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                      stop_gen();
                  else
                      re_start_gen();                      
                  continue;
              end
          end //if(nack_flag==1)
          //->i2c_if.event_master_general_call_addr_sent;
          send_byte(gen_call_second_byte);
          // check and response when addr/send_start_byte nack generated by slave    
          if(nack_flag==1) begin
              if(num_of_retry==0 | !trans.retry_if_nack) begin
                  stop_gen();
                  return;
              end
              else if(retry_num==num_of_retry) begin
                  retry_num++;
                  continue;
              end
              else begin
                  retry_num++;
                  if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                      stop_gen();
                  else
                      re_start_gen();                      
                  continue;
              end
          end
          //->i2c_if.event_master_general_call_sec_byte_sent;
          //if(gen_call_second_byte[0]==1'b1) begin
          //if send_start_byte==1,send start byte.
          
          for(int i=0; i<trans.data.size();i++)
          begin
              send_byte(trans.data[i]);
              // check and response when data nack generated by slave    
              if(nack_flag==1) begin
                  if(num_of_retry==0 | !trans.retry_if_nack) begin
                      stop_gen();
                      return;
                  end
                  else if(retry_num==num_of_retry) begin
                      retry_num++;
                      continue;
                  end
                  else begin
                      retry_num++;
                      if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                          stop_gen();
                      else
                          re_start_gen();
                      break;
                  end     
              end  //  if(nack_flag==1)           
          end
          
          if(nack_flag==0 | retry_num==num_of_retry+1) begin
              if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                  stop_gen();
              else
                  re_start_gen();
              break;
          end  //if(nack_flag==0)
      end
    I2C_DEVICE_ID: 
      for(int retry_num=0; retry_num<=num_of_retry; ) begin  
          start_gen();
          send_byte(device_id_w);
          // check and response when addr/send_start_byte nack generated by slave    
          if(nack_flag==1) begin
              if(num_of_retry==0 | !trans.retry_if_nack) begin
                  stop_gen();
                  return;
              end
              else if(retry_num==num_of_retry) begin
                  retry_num++; 
                  continue;
              end
              else begin
                  retry_num++;
                  if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                      stop_gen();
                  else
                      re_start_gen();
                  continue;
              end
          end

          if(trans.addr_10bit ==1)
              rw_slave_10bit_addr(trans.addr, 0);
          else
              rw_slave_7bit_addr(trans.addr[6:0], 0);
          //ack/noack don't care
          
          if(trans.m_device_id_gen_stop==0) begin
              re_start_gen();
              send_byte(device_id_r);
              // check and response when addr/send_start_byte nack generated by slave    
              if(nack_flag==1) begin
                  if(num_of_retry==0 | !trans.retry_if_nack) begin
                      stop_gen();
                      return;
                  end
                  else if(retry_num==num_of_retry) begin
                      retry_num++; 
                      continue;
                  end
                  else begin
                      retry_num++;
                      if(trans.sr_or_p_gen==0) //0--gen sotp, 1--gen re-start
                          stop_gen();
                      else
                          re_start_gen();
                      continue;
                  end
              end //if(nack_flag==1)

              if(trans.device_id_rollback_iteration ==0)  begin   //no rollback
                  case(trans.nack_at_device_id_byte)
                    1:
                      begin
                          recv_byte_noack(recv_data);
                          trans.data[0] = recv_data;
                          
                          if(trans.sr_or_p_gen==0  | retry_num==num_of_retry+1  | retry_num==0) begin //0--gen sotp, 1--gen re-start
                              retry_num++;
                              stop_gen();
                          end
                          else
                              re_start_gen();
                          break;                            
                      end
                    2:
                      begin
                          recv_byte(recv_data);
                          trans.data[0] = recv_data;
                          recv_byte_noack(recv_data);
                          trans.data[1] = recv_data;
                          
                          if(trans.sr_or_p_gen==0  | retry_num==num_of_retry+1  | retry_num==0) begin //0--gen sotp, 1--gen re-start
                              retry_num++;
                              stop_gen();
                          end
                          else
                              re_start_gen();
                          
                          break;
                      end
                    default:
                      begin
                          recv_byte(recv_data);
                          trans.data[0] = recv_data;
                          recv_byte(recv_data);
                          trans.data[1] = recv_data;
                          recv_byte_noack(recv_data);
                          trans.data[2] = recv_data;
                          
                          if(trans.sr_or_p_gen==0  | retry_num==num_of_retry+1  | retry_num==0) begin //0--gen sotp, 1--gen re-start
                              retry_num++;
                              stop_gen();
                          end
                          else
                              re_start_gen();
                          
                          break;
                      end
                    endcase
              end  //if(trans.device_id_rollback_iteration ==0)
              else begin    //rollback
                  for(int i=0;i<trans.nack_at_device_id_byte-1;i++) begin
                      recv_byte(recv_data);
                      trans.data[i] = recv_data;
                  end
                  recv_byte_noack(recv_data);
                  trans.data[trans.nack_at_device_id_byte-1] = recv_data;
                
                  if(trans.sr_or_p_gen==0  | retry_num==num_of_retry+1  | retry_num==0) begin //0--gen sotp, 1--gen re-start
                      retry_num++;
                      stop_gen();
                  end
                  else
                      re_start_gen();
                  
                  break;                  
              end//else begin    //rollback
          end//if(trans.m_device_id_gen_stop==0)
          else begin
              if(trans.sr_or_p_gen==0  | retry_num==num_of_retry+1  | retry_num==0) begin //0--gen sotp, 1--gen re-start
                  retry_num++;
                  stop_gen();
              end
              else
                  re_start_gen();
              break;
          end
      end
    default:  
      begin  
         `uvm_error("i2c_master_driver_common","i2c command error!!!");
      end
  endcase
endtask : drive_data

task lvc_i2c_master_driver_common::collect_response_from_vif(lvc_i2c_master_transaction trans);
  // TODO detailed bus response collection here!!!
endtask

task lvc_i2c_master_driver_common::start_gen();
  if(lock.try_get()) begin
    //repeat(1000) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 1;
    i2c_if.sda_master = 1;
    repeat(1000) @(posedge i2c_if.CLK);
    i2c_if.sda_master = 0;
    repeat(sta_hd) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 0;
    //->i2c_if.event_master_start_generated;
  end
  else 
    `uvm_info("start", "Because The Last Transaction Have Generate Restart CMD, This Transation Need Not Generate Start CMD", UVM_DEBUG);
endtask : start_gen

task lvc_i2c_master_driver_common::re_start_gen();
  //bus free time, hs mode no this parameter.
  fork
      begin
          repeat(i2c_clk_low) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
      end
      begin
          repeat(i2c_clk_low-re_sta_su) @(posedge i2c_if.CLK);
          i2c_if.sda_master = 1;
      end
  join

  repeat(re_sta_su) @(posedge i2c_if.CLK);
  i2c_if.sda_master = 0;
  repeat(sta_hd) @(posedge i2c_if.CLK);
  i2c_if.scl_master = 0;
  //->i2c_if.event_master_repeated_start_generated;
endtask : re_start_gen

task lvc_i2c_master_driver_common::pre_hs_in_fm_start_gen();
  if(lock.try_get()) begin
    repeat(cfg.scl_low_time_fs) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 1;
    i2c_if.sda_master = 1;
    repeat(cfg.scl_low_time_fs) @(posedge i2c_if.CLK);
    i2c_if.sda_master = 0;
    repeat(cfg.scl_high_time_fs) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 0;
    //->i2c_if.event_master_start_generated;
  end
  else 
    `uvm_info("start", "Because The Last Transaction Have Generate Restart CMD, This Transation Need Not Generate Start CMD", UVM_DEBUG);
endtask : pre_hs_in_fm_start_gen

task lvc_i2c_master_driver_common::pre_hs_in_fm_plus_start_gen();
  if(lock.try_get()) begin
    repeat(cfg.scl_low_time_fm_plus) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 1;
    i2c_if.sda_master = 1;
    repeat(cfg.scl_low_time_fm_plus) @(posedge i2c_if.CLK);
    i2c_if.sda_master = 0;
    repeat(cfg.scl_high_time_fm_plus) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 0;
    //->i2c_if.event_master_start_generated;
  end
  else 
    `uvm_info("start", "Because The Last Transaction Have Generate Restart CMD, This Transation Need Not Generate Start CMD", UVM_DEBUG);
endtask : pre_hs_in_fm_plus_start_gen

task lvc_i2c_master_driver_common::stop_gen();
  fork
      begin
          wait_data_hd_time();
          i2c_if.sda_master = 0;
      end
      begin
          repeat(i2c_clk_low) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
          wait(i2c_if.SCL == 1);
      end
  join
  repeat(sto_su) @(posedge i2c_if.CLK);
  i2c_if.sda_master = 1;
  repeat(tbuf_time) @(posedge i2c_if.CLK);
//  i2c_if.scl_master = 1'bz;
//  i2c_if.sda_master = 1'bz;
  //->i2c_if.event_master_stop_generated;
  lock.put();
endtask : stop_gen

task lvc_i2c_master_driver_common::rw_slave_7bit_addr(bit[6:0] addr, bit rw);
  for(int i=6;i>=0;i--) begin
    fork
      begin
          wait_data_hd_time();
          i2c_if.sda_master = addr[i];
      end
      begin
          repeat(i2c_clk_low) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
      end
    join
  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
  i2c_if.scl_master = 0;
  end
  fork
      begin
          wait_data_hd_time();
          i2c_if.sda_master = rw;
      end
      begin
          repeat(i2c_clk_low) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
      end
  join
  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
  i2c_if.scl_master = 0;
  fork
      begin
          repeat(i2c_clk_low) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
          if(i2c_if.SDA !=0)
            nack_flag = 1;
          else
            nack_flag = 0;
          //`uvm_error("master driver sent 7 bit slave addr","slave send no ack to master.")
      end
  join 
  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
  i2c_if.scl_master = 0;
endtask : rw_slave_7bit_addr

task lvc_i2c_master_driver_common::rw_slave_10bit_addr(bit [9:0] addr, bit rw);
   bit[7:0] wr_fst_byte = {5'b11110,addr[9:8],1'b0}; 
   bit[7:0] rd_fst_byte = {5'b11110,addr[9:8],1'b1}; 

   if(rw == 0)  begin  //write data to 10bits address slave
     for(int i=7;i>=0;i--) begin   //write 10bits address high 2bit
       fork
           begin
               wait_data_hd_time();
               i2c_if.sda_master = wr_fst_byte[i];
           end
           begin
               repeat(i2c_clk_low) @(posedge i2c_if.CLK);
               i2c_if.scl_master = 1;
           end
       join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     end
     fork
       begin
//         wait_data_hd_time();
//         i2c_if.sda_master = 1'bz;
       end
       begin
         repeat(i2c_clk_low) @(posedge i2c_if.CLK);
         i2c_if.scl_master = 1;
         if(i2c_if.sda_master !=0)
           nack_flag=1;
         else
           nack_flag=0;
            //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
       end
     join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);   
       i2c_if.scl_master = 0;
     
     for(int i=7;i>=0;i--) begin   //write 10bits address low 8bit
       fork
         begin
           wait_data_hd_time();
           i2c_if.sda_master = addr[i];
         end
         begin
           repeat(i2c_clk_low) @(posedge i2c_if.CLK);
           i2c_if.scl_master = 1;
         end
       join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     end
     fork
       begin
 //        wait_data_hd_time();
//         i2c_if.sda_master = 1'bz;
       end
       begin
         repeat(i2c_clk_low) @(posedge i2c_if.CLK);
         i2c_if.scl_master = 1;
         if(i2c_if.sda_master !=0)
           nack_flag=1;
         else
           nack_flag=0;
          //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
       end
     join      
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
   end 
   else begin          //read data from 10bits address slave
     for(int i=7;i>=0;i--) begin   //write 10bits address high 2bit
       fork
           begin
               wait_data_hd_time();
               i2c_if.sda_master = wr_fst_byte[i];
           end
           begin
               repeat(i2c_clk_low) @(posedge i2c_if.CLK);
               i2c_if.scl_master = 1;
           end
         join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     end
     fork
       begin
 //        wait_data_hd_time();
//         i2c_if.sda_master = 1'bz;
       end
       begin
         repeat(i2c_clk_low) @(posedge i2c_if.CLK);
         i2c_if.scl_master = 1;
         if(i2c_if.sda_master !=0)
           nack_flag=1;
         else
           nack_flag=0;
            //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
       end
     join
     repeat(i2c_clk_high) @(posedge i2c_if.CLK);
     i2c_if.scl_master = 0;
     
     for(int i=7;i>=0;i--) begin   //write 10bits address low 8bit
       fork
         begin
           wait_data_hd_time();
           i2c_if.sda_master = addr[i];
         end
         begin
           repeat(i2c_clk_low) @(posedge i2c_if.CLK);
           i2c_if.scl_master = 1;
         end
       join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     end
     fork
       begin
 //        wait_data_hd_time();
 //        i2c_if.sda_master = 1'bz;
       end
       begin
         repeat(i2c_clk_low) @(posedge i2c_if.CLK);
         i2c_if.scl_master = 1;
         if(i2c_if.sda_master !=0)
           nack_flag=1;
         else
           nack_flag=0;
            //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
        end
      join
          repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     
     re_start_gen();
     for(int i=7;i>=0;i--) begin   //write 10bits address high 2bit
       fork
         begin
           wait_data_hd_time();
           i2c_if.sda_master = rd_fst_byte[i];
         end
         begin
           repeat(i2c_clk_low) @(posedge i2c_if.CLK);
            i2c_if.scl_master = 1;
          end
        join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     end
     fork
     begin
 //      wait_data_hd_time();
 //      i2c_if.sda_master = 1'bz;
     end
     begin
       repeat(i2c_clk_low) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 1;
       if(i2c_if.sda_master !=0)
         nack_flag=1;
       else
         nack_flag=0;
          //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
        end
      join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
   end
endtask : rw_slave_10bit_addr

task lvc_i2c_master_driver_common::send_byte(bit[7:0] send_byte);
  // i2c_if.scl_master = 0;
 //  wait(i2c_if.SCL&i2c_if.SDA != 1'bz); //stretch release
  for(int i=7;i>=0;i--) begin
  fork
      begin
          wait_data_hd_time();
          i2c_if.sda_master=send_byte[i];
      end
      begin
          repeat(i2c_clk_low) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
          wait(i2c_if.SCL == 1);
      end
  join
  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
  i2c_if.scl_master = 0;
  end
  fork
      begin
 //         wait_data_hd_time();
//          i2c_if.sda_master = 1'bz;
      end
      begin
          repeat(i2c_clk_low) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
          if(i2c_if.sda_master != 0)
            nack_flag=1;
          else
            nack_flag=0;
          //`uvm_error("master driver sent byte to slave","slave send no ack to master.")
      end
  join
  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
  i2c_if.scl_master = 0;
endtask : send_byte

task lvc_i2c_master_driver_common::pre_hs_in_fm_send_byte(bit[7:0] send_byte);
  for(int i=7;i>=0;i--) begin
  fork
      begin
          repeat(cfg.min_hd_dat_time_fs) @(posedge i2c_if.CLK);
          i2c_if.sda_master=send_byte[i];
      end
      begin
          repeat(cfg.scl_low_time_fs) @(posedge i2c_if.CLK);  
          i2c_if.scl_master = 1;
      end
  join
  repeat(cfg.scl_high_time_fs) @(posedge i2c_if.CLK);  
  i2c_if.scl_master = 0;
  end
  fork
      begin
 //         repeat(cfg.min_hd_dat_time_fs) @(posedge i2c_if.CLK);
 //         i2c_if.sda_master = 1'bz;
      end
      begin
          repeat(cfg.scl_low_time_fs) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
          if(i2c_if.sda_master != 1)
          `uvm_error("master driver sent hs pre byte to slave","slave send ack to master.")
      end
  join
  repeat(cfg.scl_high_time_fs) @(posedge i2c_if.CLK);  
  i2c_if.scl_master = 0;
endtask : pre_hs_in_fm_send_byte

task lvc_i2c_master_driver_common::pre_hs_in_fm_plus_send_byte(bit[7:0] send_byte);
  for(int i=7;i>=0;i--) begin
  fork
      begin
          repeat(cfg.min_hd_dat_time_fm_plus) @(posedge i2c_if.CLK);
          i2c_if.sda_master=send_byte[i];
      end
      begin
          repeat(cfg.scl_low_time_fm_plus) @(posedge i2c_if.CLK);  
          i2c_if.scl_master = 1;
      end
  join
  repeat(cfg.scl_high_time_fm_plus) @(posedge i2c_if.CLK);  
  i2c_if.scl_master = 0;
  end
  fork
      begin
 //         repeat(cfg.min_hd_dat_time_fm_plus) @(posedge i2c_if.CLK);
 //         i2c_if.sda_master = 1'bz;
      end
      begin
          repeat(cfg.scl_low_time_fm_plus) @(posedge i2c_if.CLK);
          i2c_if.scl_master = 1;
          if(i2c_if.sda_master != 1)
          `uvm_error("master driver sent hs pre byte to slave","slave send ack to master.")
      end
  join
  repeat(cfg.scl_high_time_fm_plus) @(posedge i2c_if.CLK);  
  i2c_if.scl_master = 0;
endtask : pre_hs_in_fm_plus_send_byte

task lvc_i2c_master_driver_common::recv_byte(output bit[7:0] recv_data);
  for(int i=7;i>=0;i--) begin
    repeat(i2c_clk_low) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 1;
    // wait until the i2c slave release SCL
    wait(i2c_if.SCL === 1'b1);
    recv_data[i] = i2c_if.SDA;
    repeat(i2c_clk_high) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 0;
  end
  fork
    begin
      wait_data_hd_time();
      i2c_if.sda_master = 0;   //send ack to slave
    end
    begin
      repeat(i2c_clk_low) @(posedge i2c_if.CLK);
      i2c_if.scl_master = 1;
    end
  join
  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
  i2c_if.sda_master = 1;   // finish the data ack
  i2c_if.scl_master = 0;
endtask : recv_byte

task lvc_i2c_master_driver_common::recv_byte_noack(output bit[7:0] recv_data);  //the last data received, master will sent out a n-ack to slave
  for(int i=7;i>=0;i--) begin
    repeat(i2c_clk_low) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 1;
    recv_data[i] = i2c_if.SDA;
    repeat(i2c_clk_high) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 0;
  end
  fork
    begin
      wait_data_hd_time();
      i2c_if.sda_master = 1;   //send n-ack to slave
    end
    begin
      repeat(i2c_clk_low) @(posedge i2c_if.CLK);
      i2c_if.scl_master = 1;
    end
  join
  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
  i2c_if.scl_master = 0;
endtask : recv_byte_noack

task lvc_i2c_master_driver_common::send_start_byte();
    bit[8:0]  start_byte = 9'b000000011;
    for(int i=8;i>=0;i--) begin
      fork
          begin
              wait_data_hd_time();
              i2c_if.sda_master=start_byte[i];
          end
          begin
              repeat(i2c_clk_low) @(posedge i2c_if.CLK);
              i2c_if.scl_master = 1;
          end
      join
    repeat(i2c_clk_high) @(posedge i2c_if.CLK);
    i2c_if.scl_master = 0;
    end
    //->i2c_if.event_master_start_byte_transmited;
    re_start_gen();
endtask : send_start_byte

task lvc_i2c_master_driver_common::rw_same_slave_10bit_addr(bit [9:0] addr, bit rw);
   bit[7:0] wr_fst_byte = {5'b11110,addr[9:8],1'b0}; 
   bit[7:0] rd_fst_byte = {5'b11110,addr[9:8],1'b1}; 

   if(rw == 0)  begin  //write data to 10bits address slave
     for(int i=7;i>=0;i--) begin   //write 10bits address high 2bit
       fork
           begin
               wait_data_hd_time();
               i2c_if.sda_master = wr_fst_byte[i];
           end
           begin
               repeat(i2c_clk_low) @(posedge i2c_if.CLK);
               i2c_if.scl_master = 1;
           end
       join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     end
     fork
       begin
//         wait_data_hd_time();
//         i2c_if.sda_master = 1'bz;
       end
       begin
         repeat(i2c_clk_low) @(posedge i2c_if.CLK);
         i2c_if.scl_master = 1;
         if(i2c_if.sda_master !=0)
           nack_flag=1;
         else
           nack_flag=0;
            //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
       end
     join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);   
       i2c_if.scl_master = 0;
     
     //for(int i=7;i>=0;i--) begin   //write 10bits address low 8bit
     //  fork
     //    begin
     //      wait_data_hd_time();
     //      i2c_if.sda_master = addr[i];
     //    end
     //    begin
     //      repeat(i2c_clk_low) @(posedge i2c_if.CLK);
     //      i2c_if.scl_master = 1;
     //    end
     //  join
     //  repeat(i2c_clk_high) @(posedge i2c_if.CLK);
     //  i2c_if.scl_master = 0;
     //end
     fork
       begin
 //        wait_data_hd_time();
//         i2c_if.sda_master = 1'bz;
       end
       begin
         repeat(i2c_clk_low) @(posedge i2c_if.CLK);
         i2c_if.scl_master = 1;
         if(i2c_if.sda_master !=0)
           nack_flag=1;
         else
           nack_flag=0;
          //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
       end
     join      
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
   end 
   else begin          //read data from 10bits address slave
     for(int i=7;i>=0;i--) begin   //write 10bits address high 2bit
       fork
         begin
           wait_data_hd_time();
           i2c_if.sda_master = rd_fst_byte[i];
         end
         begin
           repeat(i2c_clk_low) @(posedge i2c_if.CLK);
            i2c_if.scl_master = 1;
          end
        join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
     end
     fork
     begin
 //      wait_data_hd_time();
 //      i2c_if.sda_master = 1'bz;
     end
     begin
       repeat(i2c_clk_low) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 1;
       if(i2c_if.sda_master !=0)
         nack_flag=1;
       else
         nack_flag=0;
          //`uvm_error("master driver sent 10 bit slave addr","slave send no ack to master.")
        end
      join
       repeat(i2c_clk_high) @(posedge i2c_if.CLK);
       i2c_if.scl_master = 0;
   end
endtask : rw_same_slave_10bit_addr

`endif // LVC_I2C_MASTER_DRIVER_COMMON_SV
